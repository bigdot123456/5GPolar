module f_calculator(
	llr_a,		// the first likelihood ratio, in fixed point
	llr_b,		// the second likelihood ratio, in fixed point
	f_result	// the likelihood ratio resulting by carrying on the f operation on the inputs
);
	input	[31:0]	first_channel;
	input	[31:0]	second_channel;
	output	[31:0]	f_result;
	
	always @ (*)
	begin
		
	end
	

endmodule
